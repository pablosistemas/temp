///////////////////////////////////////////////////////////////////////////////
// $Id: header_hash.v 3582 2008-04-10 19:53:37Z jnaous $
//
// Module: hash.v
// Project: temp 
///////////////////////////////////////////////////////////////////////////////

module hash
    #(parameter INPUT_WIDTH = 96,
      parameter OUTPUT_WIDTH = 19)
    (input [INPUT_WIDTH-1:0]       data,
     output reg [OUTPUT_WIDTH-1:0] hash_0,
     output reg [OUTPUT_WIDTH-1:0] hash_1,
     input                         clk,
     input                         reset);


////////////////////////////////////////////////////////////////////////////////
// Copyright (C) 1999-2008 Easics NV.
// This source file may be used and distributed without restriction
// provided that this copyright statement is not removed from the file
// and that any derivative work contains the original copyright notice
// and the associated disclaimer.
//
// THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
// WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
//
// Purpose : synthesizable CRC function
//   * polynomial: (0 1 3 6 7 8 10 11 13 14 16 18 19 20 22)
//   * data width: 256
//
// Info : tools@easics.be
//        http://www.easics.com
////////////////////////////////////////////////////////////////////////////////

  // polynomial: (0 1 3 6 7 8 10 11 13 14 16 18 19 20 22)
  // data width: 256
  // convention: the first serial bit is D[255]
  function [21:0] crc_func_0;

    input [255:0] Data;
    input [21:0] crc;
    reg [255:0] d;
    reg [21:0] c;
    reg [21:0] newcrc;
  begin
    d = Data;
    c = crc;

    newcrc[0] = d[255] ^ d[253] ^ d[252] ^ d[250] ^ d[249] ^ d[246] ^ d[245] ^ d[243] ^ d[242] ^ d[241] ^ d[239] ^ d[238] ^ d[237] ^ d[236] ^ d[233] ^ d[232] ^ d[228] ^ d[227] ^ d[226] ^ d[224] ^ d[222] ^ d[221] ^ d[220] ^ d[216] ^ d[215] ^ d[211] ^ d[208] ^ d[205] ^ d[204] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[199] ^ d[195] ^ d[193] ^ d[192] ^ d[191] ^ d[190] ^ d[188] ^ d[182] ^ d[181] ^ d[179] ^ d[176] ^ d[175] ^ d[174] ^ d[172] ^ d[170] ^ d[165] ^ d[162] ^ d[160] ^ d[154] ^ d[150] ^ d[148] ^ d[147] ^ d[146] ^ d[145] ^ d[143] ^ d[138] ^ d[136] ^ d[135] ^ d[128] ^ d[127] ^ d[126] ^ d[124] ^ d[123] ^ d[122] ^ d[119] ^ d[116] ^ d[114] ^ d[112] ^ d[110] ^ d[107] ^ d[106] ^ d[105] ^ d[104] ^ d[100] ^ d[99] ^ d[98] ^ d[87] ^ d[85] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[72] ^ d[71] ^ d[70] ^ d[66] ^ d[65] ^ d[63] ^ d[61] ^ d[59] ^ d[58] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[51] ^ d[50] ^ d[49] ^ d[47] ^ d[45] ^ d[44] ^ d[43] ^ d[42] ^ d[40] ^ d[39] ^ d[37] ^ d[33] ^ d[32] ^ d[31] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[16] ^ d[13] ^ d[11] ^ d[8] ^ d[7] ^ d[6] ^ d[3] ^ d[2] ^ d[0] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[7] ^ c[8] ^ c[9] ^ c[11] ^ c[12] ^ c[15] ^ c[16] ^ c[18] ^ c[19] ^ c[21];
    newcrc[1] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[249] ^ d[247] ^ d[245] ^ d[244] ^ d[241] ^ d[240] ^ d[236] ^ d[234] ^ d[232] ^ d[229] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[220] ^ d[217] ^ d[215] ^ d[212] ^ d[211] ^ d[209] ^ d[208] ^ d[206] ^ d[199] ^ d[196] ^ d[195] ^ d[194] ^ d[190] ^ d[189] ^ d[188] ^ d[183] ^ d[181] ^ d[180] ^ d[179] ^ d[177] ^ d[174] ^ d[173] ^ d[172] ^ d[171] ^ d[170] ^ d[166] ^ d[165] ^ d[163] ^ d[162] ^ d[161] ^ d[160] ^ d[155] ^ d[154] ^ d[151] ^ d[150] ^ d[149] ^ d[145] ^ d[144] ^ d[143] ^ d[139] ^ d[138] ^ d[137] ^ d[135] ^ d[129] ^ d[126] ^ d[125] ^ d[122] ^ d[120] ^ d[119] ^ d[117] ^ d[116] ^ d[115] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[110] ^ d[108] ^ d[104] ^ d[101] ^ d[98] ^ d[88] ^ d[87] ^ d[86] ^ d[85] ^ d[82] ^ d[77] ^ d[76] ^ d[75] ^ d[73] ^ d[70] ^ d[67] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[60] ^ d[58] ^ d[57] ^ d[53] ^ d[52] ^ d[49] ^ d[48] ^ d[47] ^ d[46] ^ d[42] ^ d[41] ^ d[39] ^ d[38] ^ d[37] ^ d[34] ^ d[31] ^ d[28] ^ d[18] ^ d[17] ^ d[16] ^ d[14] ^ d[13] ^ d[12] ^ d[11] ^ d[9] ^ d[6] ^ d[4] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[2] ^ c[6] ^ c[7] ^ c[10] ^ c[11] ^ c[13] ^ c[15] ^ c[17] ^ c[18] ^ c[20] ^ c[21];
    newcrc[2] = d[255] ^ d[253] ^ d[252] ^ d[250] ^ d[248] ^ d[246] ^ d[245] ^ d[242] ^ d[241] ^ d[237] ^ d[235] ^ d[233] ^ d[230] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[221] ^ d[218] ^ d[216] ^ d[213] ^ d[212] ^ d[210] ^ d[209] ^ d[207] ^ d[200] ^ d[197] ^ d[196] ^ d[195] ^ d[191] ^ d[190] ^ d[189] ^ d[184] ^ d[182] ^ d[181] ^ d[180] ^ d[178] ^ d[175] ^ d[174] ^ d[173] ^ d[172] ^ d[171] ^ d[167] ^ d[166] ^ d[164] ^ d[163] ^ d[162] ^ d[161] ^ d[156] ^ d[155] ^ d[152] ^ d[151] ^ d[150] ^ d[146] ^ d[145] ^ d[144] ^ d[140] ^ d[139] ^ d[138] ^ d[136] ^ d[130] ^ d[127] ^ d[126] ^ d[123] ^ d[121] ^ d[120] ^ d[118] ^ d[117] ^ d[116] ^ d[115] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[109] ^ d[105] ^ d[102] ^ d[99] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[83] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[71] ^ d[68] ^ d[66] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[59] ^ d[58] ^ d[54] ^ d[53] ^ d[50] ^ d[49] ^ d[48] ^ d[47] ^ d[43] ^ d[42] ^ d[40] ^ d[39] ^ d[38] ^ d[35] ^ d[32] ^ d[29] ^ d[19] ^ d[18] ^ d[17] ^ d[15] ^ d[14] ^ d[13] ^ d[12] ^ d[10] ^ d[7] ^ d[5] ^ d[3] ^ d[2] ^ d[1] ^ c[1] ^ c[3] ^ c[7] ^ c[8] ^ c[11] ^ c[12] ^ c[14] ^ c[16] ^ c[18] ^ c[19] ^ c[21];
    newcrc[3] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[250] ^ d[247] ^ d[245] ^ d[241] ^ d[239] ^ d[237] ^ d[234] ^ d[233] ^ d[232] ^ d[231] ^ d[225] ^ d[224] ^ d[221] ^ d[220] ^ d[219] ^ d[217] ^ d[216] ^ d[215] ^ d[214] ^ d[213] ^ d[210] ^ d[205] ^ d[204] ^ d[203] ^ d[202] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[196] ^ d[195] ^ d[193] ^ d[188] ^ d[185] ^ d[183] ^ d[173] ^ d[170] ^ d[168] ^ d[167] ^ d[164] ^ d[163] ^ d[160] ^ d[157] ^ d[156] ^ d[154] ^ d[153] ^ d[152] ^ d[151] ^ d[150] ^ d[148] ^ d[143] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[136] ^ d[135] ^ d[131] ^ d[126] ^ d[123] ^ d[121] ^ d[118] ^ d[117] ^ d[115] ^ d[113] ^ d[107] ^ d[105] ^ d[104] ^ d[103] ^ d[99] ^ d[98] ^ d[90] ^ d[89] ^ d[88] ^ d[85] ^ d[84] ^ d[81] ^ d[80] ^ d[71] ^ d[70] ^ d[69] ^ d[67] ^ d[64] ^ d[62] ^ d[61] ^ d[60] ^ d[58] ^ d[56] ^ d[53] ^ d[48] ^ d[47] ^ d[45] ^ d[42] ^ d[41] ^ d[37] ^ d[36] ^ d[32] ^ d[31] ^ d[30] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[15] ^ d[14] ^ d[7] ^ d[4] ^ d[0] ^ c[0] ^ c[3] ^ c[5] ^ c[7] ^ c[11] ^ c[13] ^ c[16] ^ c[17] ^ c[18] ^ c[20] ^ c[21];
    newcrc[4] = d[255] ^ d[253] ^ d[252] ^ d[251] ^ d[248] ^ d[246] ^ d[242] ^ d[240] ^ d[238] ^ d[235] ^ d[234] ^ d[233] ^ d[232] ^ d[226] ^ d[225] ^ d[222] ^ d[221] ^ d[220] ^ d[218] ^ d[217] ^ d[216] ^ d[215] ^ d[214] ^ d[211] ^ d[206] ^ d[205] ^ d[204] ^ d[203] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[196] ^ d[194] ^ d[189] ^ d[186] ^ d[184] ^ d[174] ^ d[171] ^ d[169] ^ d[168] ^ d[165] ^ d[164] ^ d[161] ^ d[158] ^ d[157] ^ d[155] ^ d[154] ^ d[153] ^ d[152] ^ d[151] ^ d[149] ^ d[144] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[136] ^ d[132] ^ d[127] ^ d[124] ^ d[122] ^ d[119] ^ d[118] ^ d[116] ^ d[114] ^ d[108] ^ d[106] ^ d[105] ^ d[104] ^ d[100] ^ d[99] ^ d[91] ^ d[90] ^ d[89] ^ d[86] ^ d[85] ^ d[82] ^ d[81] ^ d[72] ^ d[71] ^ d[70] ^ d[68] ^ d[65] ^ d[63] ^ d[62] ^ d[61] ^ d[59] ^ d[57] ^ d[54] ^ d[49] ^ d[48] ^ d[46] ^ d[43] ^ d[42] ^ d[38] ^ d[37] ^ d[33] ^ d[32] ^ d[31] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[16] ^ d[15] ^ d[8] ^ d[5] ^ d[1] ^ c[0] ^ c[1] ^ c[4] ^ c[6] ^ c[8] ^ c[12] ^ c[14] ^ c[17] ^ c[18] ^ c[19] ^ c[21];
    newcrc[5] = d[254] ^ d[253] ^ d[252] ^ d[249] ^ d[247] ^ d[243] ^ d[241] ^ d[239] ^ d[236] ^ d[235] ^ d[234] ^ d[233] ^ d[227] ^ d[226] ^ d[223] ^ d[222] ^ d[221] ^ d[219] ^ d[218] ^ d[217] ^ d[216] ^ d[215] ^ d[212] ^ d[207] ^ d[206] ^ d[205] ^ d[204] ^ d[202] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[195] ^ d[190] ^ d[187] ^ d[185] ^ d[175] ^ d[172] ^ d[170] ^ d[169] ^ d[166] ^ d[165] ^ d[162] ^ d[159] ^ d[158] ^ d[156] ^ d[155] ^ d[154] ^ d[153] ^ d[152] ^ d[150] ^ d[145] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[133] ^ d[128] ^ d[125] ^ d[123] ^ d[120] ^ d[119] ^ d[117] ^ d[115] ^ d[109] ^ d[107] ^ d[106] ^ d[105] ^ d[101] ^ d[100] ^ d[92] ^ d[91] ^ d[90] ^ d[87] ^ d[86] ^ d[83] ^ d[82] ^ d[73] ^ d[72] ^ d[71] ^ d[69] ^ d[66] ^ d[64] ^ d[63] ^ d[62] ^ d[60] ^ d[58] ^ d[55] ^ d[50] ^ d[49] ^ d[47] ^ d[44] ^ d[43] ^ d[39] ^ d[38] ^ d[34] ^ d[33] ^ d[32] ^ d[29] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[17] ^ d[16] ^ d[9] ^ d[6] ^ d[2] ^ c[0] ^ c[1] ^ c[2] ^ c[5] ^ c[7] ^ c[9] ^ c[13] ^ c[15] ^ c[18] ^ c[19] ^ c[20];
    newcrc[6] = d[254] ^ d[252] ^ d[249] ^ d[248] ^ d[246] ^ d[245] ^ d[244] ^ d[243] ^ d[241] ^ d[240] ^ d[239] ^ d[238] ^ d[235] ^ d[234] ^ d[233] ^ d[232] ^ d[226] ^ d[223] ^ d[221] ^ d[219] ^ d[218] ^ d[217] ^ d[215] ^ d[213] ^ d[211] ^ d[207] ^ d[206] ^ d[204] ^ d[198] ^ d[196] ^ d[195] ^ d[193] ^ d[192] ^ d[190] ^ d[186] ^ d[182] ^ d[181] ^ d[179] ^ d[175] ^ d[174] ^ d[173] ^ d[172] ^ d[171] ^ d[167] ^ d[166] ^ d[165] ^ d[163] ^ d[162] ^ d[159] ^ d[157] ^ d[156] ^ d[155] ^ d[153] ^ d[151] ^ d[150] ^ d[148] ^ d[147] ^ d[145] ^ d[144] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[136] ^ d[135] ^ d[134] ^ d[129] ^ d[128] ^ d[127] ^ d[123] ^ d[122] ^ d[121] ^ d[120] ^ d[119] ^ d[118] ^ d[114] ^ d[112] ^ d[108] ^ d[105] ^ d[104] ^ d[102] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[93] ^ d[92] ^ d[91] ^ d[88] ^ d[85] ^ d[84] ^ d[83] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[74] ^ d[73] ^ d[71] ^ d[67] ^ d[66] ^ d[64] ^ d[58] ^ d[55] ^ d[54] ^ d[53] ^ d[49] ^ d[48] ^ d[47] ^ d[43] ^ d[42] ^ d[37] ^ d[35] ^ d[34] ^ d[32] ^ d[31] ^ d[30] ^ d[29] ^ d[28] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[17] ^ d[16] ^ d[13] ^ d[11] ^ d[10] ^ d[8] ^ d[6] ^ d[2] ^ d[0] ^ c[0] ^ c[1] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[14] ^ c[15] ^ c[18] ^ c[20];
    newcrc[7] = d[252] ^ d[247] ^ d[244] ^ d[243] ^ d[240] ^ d[238] ^ d[237] ^ d[235] ^ d[234] ^ d[232] ^ d[228] ^ d[226] ^ d[221] ^ d[219] ^ d[218] ^ d[215] ^ d[214] ^ d[212] ^ d[211] ^ d[207] ^ d[204] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[197] ^ d[196] ^ d[195] ^ d[194] ^ d[192] ^ d[190] ^ d[188] ^ d[187] ^ d[183] ^ d[181] ^ d[180] ^ d[179] ^ d[173] ^ d[170] ^ d[168] ^ d[167] ^ d[166] ^ d[165] ^ d[164] ^ d[163] ^ d[162] ^ d[158] ^ d[157] ^ d[156] ^ d[152] ^ d[151] ^ d[150] ^ d[149] ^ d[147] ^ d[142] ^ d[141] ^ d[140] ^ d[138] ^ d[137] ^ d[130] ^ d[129] ^ d[127] ^ d[126] ^ d[121] ^ d[120] ^ d[116] ^ d[115] ^ d[114] ^ d[113] ^ d[112] ^ d[110] ^ d[109] ^ d[107] ^ d[104] ^ d[103] ^ d[102] ^ d[101] ^ d[98] ^ d[94] ^ d[93] ^ d[92] ^ d[89] ^ d[87] ^ d[86] ^ d[84] ^ d[82] ^ d[77] ^ d[76] ^ d[74] ^ d[71] ^ d[70] ^ d[68] ^ d[67] ^ d[66] ^ d[63] ^ d[61] ^ d[58] ^ d[53] ^ d[51] ^ d[48] ^ d[47] ^ d[45] ^ d[42] ^ d[40] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[30] ^ d[29] ^ d[27] ^ d[26] ^ d[25] ^ d[19] ^ d[17] ^ d[16] ^ d[14] ^ d[13] ^ d[12] ^ d[9] ^ d[8] ^ d[6] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[3] ^ c[4] ^ c[6] ^ c[9] ^ c[10] ^ c[13] ^ c[18];
    newcrc[8] = d[255] ^ d[252] ^ d[250] ^ d[249] ^ d[248] ^ d[246] ^ d[244] ^ d[243] ^ d[242] ^ d[237] ^ d[235] ^ d[232] ^ d[229] ^ d[228] ^ d[226] ^ d[224] ^ d[221] ^ d[219] ^ d[213] ^ d[212] ^ d[211] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[196] ^ d[192] ^ d[190] ^ d[189] ^ d[184] ^ d[180] ^ d[179] ^ d[176] ^ d[175] ^ d[172] ^ d[171] ^ d[170] ^ d[169] ^ d[168] ^ d[167] ^ d[166] ^ d[164] ^ d[163] ^ d[162] ^ d[160] ^ d[159] ^ d[158] ^ d[157] ^ d[154] ^ d[153] ^ d[152] ^ d[151] ^ d[147] ^ d[146] ^ d[145] ^ d[142] ^ d[141] ^ d[139] ^ d[136] ^ d[135] ^ d[131] ^ d[130] ^ d[126] ^ d[124] ^ d[123] ^ d[121] ^ d[119] ^ d[117] ^ d[115] ^ d[113] ^ d[112] ^ d[111] ^ d[108] ^ d[107] ^ d[106] ^ d[103] ^ d[102] ^ d[100] ^ d[98] ^ d[95] ^ d[94] ^ d[93] ^ d[90] ^ d[88] ^ d[83] ^ d[81] ^ d[80] ^ d[79] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[58] ^ d[56] ^ d[55] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[45] ^ d[44] ^ d[42] ^ d[41] ^ d[38] ^ d[36] ^ d[33] ^ d[32] ^ d[30] ^ d[28] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[19] ^ d[17] ^ d[16] ^ d[15] ^ d[14] ^ d[11] ^ d[10] ^ d[9] ^ d[8] ^ d[6] ^ d[1] ^ d[0] ^ c[1] ^ c[3] ^ c[8] ^ c[9] ^ c[10] ^ c[12] ^ c[14] ^ c[15] ^ c[16] ^ c[18] ^ c[21];
    newcrc[9] = d[253] ^ d[251] ^ d[250] ^ d[249] ^ d[247] ^ d[245] ^ d[244] ^ d[243] ^ d[238] ^ d[236] ^ d[233] ^ d[230] ^ d[229] ^ d[227] ^ d[225] ^ d[222] ^ d[220] ^ d[214] ^ d[213] ^ d[212] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[193] ^ d[191] ^ d[190] ^ d[185] ^ d[181] ^ d[180] ^ d[177] ^ d[176] ^ d[173] ^ d[172] ^ d[171] ^ d[170] ^ d[169] ^ d[168] ^ d[167] ^ d[165] ^ d[164] ^ d[163] ^ d[161] ^ d[160] ^ d[159] ^ d[158] ^ d[155] ^ d[154] ^ d[153] ^ d[152] ^ d[148] ^ d[147] ^ d[146] ^ d[143] ^ d[142] ^ d[140] ^ d[137] ^ d[136] ^ d[132] ^ d[131] ^ d[127] ^ d[125] ^ d[124] ^ d[122] ^ d[120] ^ d[118] ^ d[116] ^ d[114] ^ d[113] ^ d[112] ^ d[109] ^ d[108] ^ d[107] ^ d[104] ^ d[103] ^ d[101] ^ d[99] ^ d[96] ^ d[95] ^ d[94] ^ d[91] ^ d[89] ^ d[84] ^ d[82] ^ d[81] ^ d[80] ^ d[71] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[59] ^ d[57] ^ d[56] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[49] ^ d[48] ^ d[47] ^ d[46] ^ d[45] ^ d[43] ^ d[42] ^ d[39] ^ d[37] ^ d[34] ^ d[33] ^ d[31] ^ d[29] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[20] ^ d[18] ^ d[17] ^ d[16] ^ d[15] ^ d[12] ^ d[11] ^ d[10] ^ d[9] ^ d[7] ^ d[2] ^ d[1] ^ c[2] ^ c[4] ^ c[9] ^ c[10] ^ c[11] ^ c[13] ^ c[15] ^ c[16] ^ c[17] ^ c[19];
    newcrc[10] = d[255] ^ d[254] ^ d[253] ^ d[251] ^ d[249] ^ d[248] ^ d[244] ^ d[243] ^ d[242] ^ d[241] ^ d[238] ^ d[236] ^ d[234] ^ d[233] ^ d[232] ^ d[231] ^ d[230] ^ d[227] ^ d[224] ^ d[223] ^ d[222] ^ d[220] ^ d[216] ^ d[214] ^ d[213] ^ d[211] ^ d[208] ^ d[205] ^ d[204] ^ d[203] ^ d[198] ^ d[195] ^ d[194] ^ d[193] ^ d[190] ^ d[188] ^ d[186] ^ d[179] ^ d[178] ^ d[177] ^ d[176] ^ d[175] ^ d[173] ^ d[171] ^ d[169] ^ d[168] ^ d[166] ^ d[164] ^ d[161] ^ d[159] ^ d[156] ^ d[155] ^ d[153] ^ d[150] ^ d[149] ^ d[146] ^ d[145] ^ d[144] ^ d[141] ^ d[137] ^ d[136] ^ d[135] ^ d[133] ^ d[132] ^ d[127] ^ d[125] ^ d[124] ^ d[122] ^ d[121] ^ d[117] ^ d[116] ^ d[115] ^ d[113] ^ d[112] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[102] ^ d[99] ^ d[98] ^ d[97] ^ d[96] ^ d[95] ^ d[92] ^ d[90] ^ d[87] ^ d[83] ^ d[82] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[69] ^ d[68] ^ d[67] ^ d[64] ^ d[61] ^ d[60] ^ d[59] ^ d[57] ^ d[56] ^ d[52] ^ d[51] ^ d[48] ^ d[46] ^ d[45] ^ d[42] ^ d[39] ^ d[38] ^ d[37] ^ d[35] ^ d[34] ^ d[33] ^ d[31] ^ d[30] ^ d[22] ^ d[20] ^ d[17] ^ d[12] ^ d[10] ^ d[7] ^ d[6] ^ d[0] ^ c[0] ^ c[2] ^ c[4] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[14] ^ c[15] ^ c[17] ^ c[19] ^ c[20] ^ c[21];
    newcrc[11] = d[254] ^ d[253] ^ d[246] ^ d[244] ^ d[241] ^ d[238] ^ d[236] ^ d[235] ^ d[234] ^ d[231] ^ d[227] ^ d[226] ^ d[225] ^ d[223] ^ d[222] ^ d[220] ^ d[217] ^ d[216] ^ d[214] ^ d[212] ^ d[211] ^ d[209] ^ d[208] ^ d[206] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[196] ^ d[194] ^ d[193] ^ d[192] ^ d[190] ^ d[189] ^ d[188] ^ d[187] ^ d[182] ^ d[181] ^ d[180] ^ d[178] ^ d[177] ^ d[175] ^ d[169] ^ d[167] ^ d[157] ^ d[156] ^ d[151] ^ d[148] ^ d[143] ^ d[142] ^ d[137] ^ d[135] ^ d[134] ^ d[133] ^ d[127] ^ d[125] ^ d[124] ^ d[119] ^ d[118] ^ d[117] ^ d[113] ^ d[112] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[104] ^ d[103] ^ d[97] ^ d[96] ^ d[93] ^ d[91] ^ d[88] ^ d[87] ^ d[85] ^ d[84] ^ d[83] ^ d[77] ^ d[76] ^ d[75] ^ d[72] ^ d[71] ^ d[69] ^ d[68] ^ d[66] ^ d[63] ^ d[62] ^ d[60] ^ d[59] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[46] ^ d[45] ^ d[44] ^ d[42] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[34] ^ d[33] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[22] ^ d[20] ^ d[19] ^ d[16] ^ d[6] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[4] ^ c[7] ^ c[10] ^ c[12] ^ c[19] ^ c[20];
    newcrc[12] = d[255] ^ d[254] ^ d[247] ^ d[245] ^ d[242] ^ d[239] ^ d[237] ^ d[236] ^ d[235] ^ d[232] ^ d[228] ^ d[227] ^ d[226] ^ d[224] ^ d[223] ^ d[221] ^ d[218] ^ d[217] ^ d[215] ^ d[213] ^ d[212] ^ d[210] ^ d[209] ^ d[207] ^ d[204] ^ d[203] ^ d[202] ^ d[201] ^ d[197] ^ d[195] ^ d[194] ^ d[193] ^ d[191] ^ d[190] ^ d[189] ^ d[188] ^ d[183] ^ d[182] ^ d[181] ^ d[179] ^ d[178] ^ d[176] ^ d[170] ^ d[168] ^ d[158] ^ d[157] ^ d[152] ^ d[149] ^ d[144] ^ d[143] ^ d[138] ^ d[136] ^ d[135] ^ d[134] ^ d[128] ^ d[126] ^ d[125] ^ d[120] ^ d[119] ^ d[118] ^ d[114] ^ d[113] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[105] ^ d[104] ^ d[98] ^ d[97] ^ d[94] ^ d[92] ^ d[89] ^ d[88] ^ d[86] ^ d[85] ^ d[84] ^ d[78] ^ d[77] ^ d[76] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[67] ^ d[64] ^ d[63] ^ d[61] ^ d[60] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[53] ^ d[52] ^ d[51] ^ d[47] ^ d[46] ^ d[45] ^ d[43] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[34] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[23] ^ d[21] ^ d[20] ^ d[17] ^ d[7] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ c[1] ^ c[2] ^ c[3] ^ c[5] ^ c[8] ^ c[11] ^ c[13] ^ c[20] ^ c[21];
    newcrc[13] = d[253] ^ d[252] ^ d[250] ^ d[249] ^ d[248] ^ d[245] ^ d[242] ^ d[241] ^ d[240] ^ d[239] ^ d[232] ^ d[229] ^ d[226] ^ d[225] ^ d[221] ^ d[220] ^ d[219] ^ d[218] ^ d[215] ^ d[214] ^ d[213] ^ d[210] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[196] ^ d[194] ^ d[193] ^ d[189] ^ d[188] ^ d[184] ^ d[183] ^ d[181] ^ d[180] ^ d[177] ^ d[176] ^ d[175] ^ d[174] ^ d[172] ^ d[171] ^ d[170] ^ d[169] ^ d[165] ^ d[162] ^ d[160] ^ d[159] ^ d[158] ^ d[154] ^ d[153] ^ d[148] ^ d[147] ^ d[146] ^ d[144] ^ d[143] ^ d[139] ^ d[138] ^ d[137] ^ d[129] ^ d[128] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[120] ^ d[116] ^ d[115] ^ d[112] ^ d[111] ^ d[108] ^ d[104] ^ d[100] ^ d[95] ^ d[93] ^ d[90] ^ d[89] ^ d[86] ^ d[81] ^ d[80] ^ d[75] ^ d[74] ^ d[73] ^ d[72] ^ d[68] ^ d[66] ^ d[64] ^ d[63] ^ d[62] ^ d[57] ^ d[55] ^ d[52] ^ d[51] ^ d[50] ^ d[49] ^ d[48] ^ d[46] ^ d[45] ^ d[43] ^ d[42] ^ d[38] ^ d[36] ^ d[35] ^ d[33] ^ d[32] ^ d[31] ^ d[29] ^ d[28] ^ d[25] ^ d[23] ^ d[20] ^ d[19] ^ d[16] ^ d[13] ^ d[11] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[0] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[11] ^ c[14] ^ c[15] ^ c[16] ^ c[18] ^ c[19];
    newcrc[14] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[245] ^ d[240] ^ d[239] ^ d[238] ^ d[237] ^ d[236] ^ d[232] ^ d[230] ^ d[228] ^ d[224] ^ d[219] ^ d[214] ^ d[208] ^ d[205] ^ d[204] ^ d[203] ^ d[197] ^ d[194] ^ d[193] ^ d[192] ^ d[191] ^ d[189] ^ d[188] ^ d[185] ^ d[184] ^ d[179] ^ d[178] ^ d[177] ^ d[174] ^ d[173] ^ d[171] ^ d[166] ^ d[165] ^ d[163] ^ d[162] ^ d[161] ^ d[159] ^ d[155] ^ d[150] ^ d[149] ^ d[146] ^ d[144] ^ d[143] ^ d[140] ^ d[139] ^ d[136] ^ d[135] ^ d[130] ^ d[129] ^ d[128] ^ d[127] ^ d[126] ^ d[125] ^ d[121] ^ d[119] ^ d[117] ^ d[114] ^ d[113] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[104] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[96] ^ d[94] ^ d[91] ^ d[90] ^ d[85] ^ d[82] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[73] ^ d[72] ^ d[71] ^ d[70] ^ d[69] ^ d[67] ^ d[66] ^ d[64] ^ d[61] ^ d[59] ^ d[55] ^ d[54] ^ d[52] ^ d[46] ^ d[45] ^ d[42] ^ d[40] ^ d[36] ^ d[34] ^ d[31] ^ d[30] ^ d[29] ^ d[27] ^ d[25] ^ d[23] ^ d[22] ^ d[19] ^ d[18] ^ d[17] ^ d[16] ^ d[14] ^ d[13] ^ d[12] ^ d[11] ^ d[5] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[11] ^ c[17] ^ c[18] ^ c[20] ^ c[21];
    newcrc[15] = d[255] ^ d[253] ^ d[252] ^ d[246] ^ d[241] ^ d[240] ^ d[239] ^ d[238] ^ d[237] ^ d[233] ^ d[231] ^ d[229] ^ d[225] ^ d[220] ^ d[215] ^ d[209] ^ d[206] ^ d[205] ^ d[204] ^ d[198] ^ d[195] ^ d[194] ^ d[193] ^ d[192] ^ d[190] ^ d[189] ^ d[186] ^ d[185] ^ d[180] ^ d[179] ^ d[178] ^ d[175] ^ d[174] ^ d[172] ^ d[167] ^ d[166] ^ d[164] ^ d[163] ^ d[162] ^ d[160] ^ d[156] ^ d[151] ^ d[150] ^ d[147] ^ d[145] ^ d[144] ^ d[141] ^ d[140] ^ d[137] ^ d[136] ^ d[131] ^ d[130] ^ d[129] ^ d[128] ^ d[127] ^ d[126] ^ d[122] ^ d[120] ^ d[118] ^ d[115] ^ d[114] ^ d[111] ^ d[110] ^ d[108] ^ d[107] ^ d[105] ^ d[102] ^ d[101] ^ d[100] ^ d[99] ^ d[97] ^ d[95] ^ d[92] ^ d[91] ^ d[86] ^ d[83] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[74] ^ d[73] ^ d[72] ^ d[71] ^ d[70] ^ d[68] ^ d[67] ^ d[65] ^ d[62] ^ d[60] ^ d[56] ^ d[55] ^ d[53] ^ d[47] ^ d[46] ^ d[43] ^ d[41] ^ d[37] ^ d[35] ^ d[32] ^ d[31] ^ d[30] ^ d[28] ^ d[26] ^ d[24] ^ d[23] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[15] ^ d[14] ^ d[13] ^ d[12] ^ d[6] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[12] ^ c[18] ^ c[19] ^ c[21];
    newcrc[16] = d[255] ^ d[254] ^ d[252] ^ d[250] ^ d[249] ^ d[247] ^ d[246] ^ d[245] ^ d[243] ^ d[240] ^ d[237] ^ d[236] ^ d[234] ^ d[233] ^ d[230] ^ d[228] ^ d[227] ^ d[224] ^ d[222] ^ d[220] ^ d[215] ^ d[211] ^ d[210] ^ d[208] ^ d[207] ^ d[206] ^ d[204] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[196] ^ d[194] ^ d[192] ^ d[188] ^ d[187] ^ d[186] ^ d[182] ^ d[180] ^ d[174] ^ d[173] ^ d[172] ^ d[170] ^ d[168] ^ d[167] ^ d[164] ^ d[163] ^ d[162] ^ d[161] ^ d[160] ^ d[157] ^ d[154] ^ d[152] ^ d[151] ^ d[150] ^ d[147] ^ d[143] ^ d[142] ^ d[141] ^ d[137] ^ d[136] ^ d[135] ^ d[132] ^ d[131] ^ d[130] ^ d[129] ^ d[126] ^ d[124] ^ d[122] ^ d[121] ^ d[115] ^ d[114] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[103] ^ d[102] ^ d[101] ^ d[99] ^ d[96] ^ d[93] ^ d[92] ^ d[85] ^ d[84] ^ d[82] ^ d[77] ^ d[76] ^ d[74] ^ d[73] ^ d[70] ^ d[69] ^ d[68] ^ d[65] ^ d[59] ^ d[58] ^ d[57] ^ d[55] ^ d[53] ^ d[51] ^ d[50] ^ d[49] ^ d[48] ^ d[45] ^ d[43] ^ d[40] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[29] ^ d[26] ^ d[23] ^ d[22] ^ d[15] ^ d[14] ^ d[11] ^ d[8] ^ d[6] ^ d[5] ^ d[4] ^ d[0] ^ c[0] ^ c[2] ^ c[3] ^ c[6] ^ c[9] ^ c[11] ^ c[12] ^ c[13] ^ c[15] ^ c[16] ^ c[18] ^ c[20] ^ c[21];
    newcrc[17] = d[255] ^ d[253] ^ d[251] ^ d[250] ^ d[248] ^ d[247] ^ d[246] ^ d[244] ^ d[241] ^ d[238] ^ d[237] ^ d[235] ^ d[234] ^ d[231] ^ d[229] ^ d[228] ^ d[225] ^ d[223] ^ d[221] ^ d[216] ^ d[212] ^ d[211] ^ d[209] ^ d[208] ^ d[207] ^ d[205] ^ d[204] ^ d[203] ^ d[202] ^ d[201] ^ d[197] ^ d[195] ^ d[193] ^ d[189] ^ d[188] ^ d[187] ^ d[183] ^ d[181] ^ d[175] ^ d[174] ^ d[173] ^ d[171] ^ d[169] ^ d[168] ^ d[165] ^ d[164] ^ d[163] ^ d[162] ^ d[161] ^ d[158] ^ d[155] ^ d[153] ^ d[152] ^ d[151] ^ d[148] ^ d[144] ^ d[143] ^ d[142] ^ d[138] ^ d[137] ^ d[136] ^ d[133] ^ d[132] ^ d[131] ^ d[130] ^ d[127] ^ d[125] ^ d[123] ^ d[122] ^ d[116] ^ d[115] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[104] ^ d[103] ^ d[102] ^ d[100] ^ d[97] ^ d[94] ^ d[93] ^ d[86] ^ d[85] ^ d[83] ^ d[78] ^ d[77] ^ d[75] ^ d[74] ^ d[71] ^ d[70] ^ d[69] ^ d[66] ^ d[60] ^ d[59] ^ d[58] ^ d[56] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[49] ^ d[46] ^ d[44] ^ d[41] ^ d[40] ^ d[39] ^ d[38] ^ d[37] ^ d[30] ^ d[27] ^ d[24] ^ d[23] ^ d[16] ^ d[15] ^ d[12] ^ d[9] ^ d[7] ^ d[6] ^ d[5] ^ d[1] ^ c[0] ^ c[1] ^ c[3] ^ c[4] ^ c[7] ^ c[10] ^ c[12] ^ c[13] ^ c[14] ^ c[16] ^ c[17] ^ c[19] ^ c[21];
    newcrc[18] = d[255] ^ d[254] ^ d[253] ^ d[251] ^ d[250] ^ d[248] ^ d[247] ^ d[246] ^ d[243] ^ d[241] ^ d[237] ^ d[235] ^ d[233] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[221] ^ d[220] ^ d[217] ^ d[216] ^ d[215] ^ d[213] ^ d[212] ^ d[211] ^ d[210] ^ d[209] ^ d[206] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[196] ^ d[195] ^ d[194] ^ d[193] ^ d[192] ^ d[191] ^ d[189] ^ d[184] ^ d[181] ^ d[179] ^ d[169] ^ d[166] ^ d[164] ^ d[163] ^ d[160] ^ d[159] ^ d[156] ^ d[153] ^ d[152] ^ d[150] ^ d[149] ^ d[148] ^ d[147] ^ d[146] ^ d[144] ^ d[139] ^ d[137] ^ d[136] ^ d[135] ^ d[134] ^ d[133] ^ d[132] ^ d[131] ^ d[127] ^ d[122] ^ d[119] ^ d[117] ^ d[114] ^ d[113] ^ d[111] ^ d[109] ^ d[103] ^ d[101] ^ d[100] ^ d[99] ^ d[95] ^ d[94] ^ d[86] ^ d[85] ^ d[84] ^ d[81] ^ d[80] ^ d[77] ^ d[76] ^ d[67] ^ d[66] ^ d[65] ^ d[63] ^ d[60] ^ d[58] ^ d[57] ^ d[56] ^ d[54] ^ d[52] ^ d[49] ^ d[44] ^ d[43] ^ d[41] ^ d[38] ^ d[37] ^ d[33] ^ d[32] ^ d[28] ^ d[27] ^ d[26] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[11] ^ d[10] ^ d[3] ^ d[0] ^ c[1] ^ c[3] ^ c[7] ^ c[9] ^ c[12] ^ c[13] ^ c[14] ^ c[16] ^ c[17] ^ c[19] ^ c[20] ^ c[21];
    newcrc[19] = d[254] ^ d[253] ^ d[251] ^ d[250] ^ d[248] ^ d[247] ^ d[246] ^ d[245] ^ d[244] ^ d[243] ^ d[241] ^ d[239] ^ d[237] ^ d[234] ^ d[233] ^ d[232] ^ d[231] ^ d[230] ^ d[229] ^ d[227] ^ d[226] ^ d[224] ^ d[220] ^ d[218] ^ d[217] ^ d[215] ^ d[214] ^ d[213] ^ d[212] ^ d[210] ^ d[208] ^ d[207] ^ d[205] ^ d[204] ^ d[203] ^ d[197] ^ d[196] ^ d[194] ^ d[191] ^ d[188] ^ d[185] ^ d[181] ^ d[180] ^ d[179] ^ d[176] ^ d[175] ^ d[174] ^ d[172] ^ d[167] ^ d[164] ^ d[162] ^ d[161] ^ d[157] ^ d[153] ^ d[151] ^ d[149] ^ d[146] ^ d[143] ^ d[140] ^ d[137] ^ d[134] ^ d[133] ^ d[132] ^ d[127] ^ d[126] ^ d[124] ^ d[122] ^ d[120] ^ d[119] ^ d[118] ^ d[116] ^ d[115] ^ d[107] ^ d[106] ^ d[105] ^ d[102] ^ d[101] ^ d[99] ^ d[98] ^ d[96] ^ d[95] ^ d[86] ^ d[82] ^ d[80] ^ d[79] ^ d[75] ^ d[72] ^ d[71] ^ d[70] ^ d[68] ^ d[67] ^ d[65] ^ d[64] ^ d[63] ^ d[57] ^ d[56] ^ d[54] ^ d[51] ^ d[49] ^ d[47] ^ d[43] ^ d[40] ^ d[38] ^ d[37] ^ d[34] ^ d[32] ^ d[31] ^ d[29] ^ d[28] ^ d[26] ^ d[25] ^ d[16] ^ d[13] ^ d[12] ^ d[8] ^ d[7] ^ d[6] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[3] ^ c[5] ^ c[7] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[16] ^ c[17] ^ c[19] ^ c[20];
    newcrc[20] = d[254] ^ d[253] ^ d[251] ^ d[250] ^ d[248] ^ d[247] ^ d[244] ^ d[243] ^ d[241] ^ d[240] ^ d[239] ^ d[237] ^ d[236] ^ d[235] ^ d[234] ^ d[231] ^ d[230] ^ d[226] ^ d[225] ^ d[224] ^ d[222] ^ d[220] ^ d[219] ^ d[218] ^ d[214] ^ d[213] ^ d[209] ^ d[206] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[193] ^ d[191] ^ d[190] ^ d[189] ^ d[188] ^ d[186] ^ d[180] ^ d[179] ^ d[177] ^ d[174] ^ d[173] ^ d[172] ^ d[170] ^ d[168] ^ d[163] ^ d[160] ^ d[158] ^ d[152] ^ d[148] ^ d[146] ^ d[145] ^ d[144] ^ d[143] ^ d[141] ^ d[136] ^ d[134] ^ d[133] ^ d[126] ^ d[125] ^ d[124] ^ d[122] ^ d[121] ^ d[120] ^ d[117] ^ d[114] ^ d[112] ^ d[110] ^ d[108] ^ d[105] ^ d[104] ^ d[103] ^ d[102] ^ d[98] ^ d[97] ^ d[96] ^ d[85] ^ d[83] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[75] ^ d[73] ^ d[70] ^ d[69] ^ d[68] ^ d[64] ^ d[63] ^ d[61] ^ d[59] ^ d[57] ^ d[56] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[49] ^ d[48] ^ d[47] ^ d[45] ^ d[43] ^ d[42] ^ d[41] ^ d[40] ^ d[38] ^ d[37] ^ d[35] ^ d[31] ^ d[30] ^ d[29] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[16] ^ d[14] ^ d[11] ^ d[9] ^ d[6] ^ d[5] ^ d[4] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[5] ^ c[6] ^ c[7] ^ c[9] ^ c[10] ^ c[13] ^ c[14] ^ c[16] ^ c[17] ^ c[19] ^ c[20];
    newcrc[21] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[249] ^ d[248] ^ d[245] ^ d[244] ^ d[242] ^ d[241] ^ d[240] ^ d[238] ^ d[237] ^ d[236] ^ d[235] ^ d[232] ^ d[231] ^ d[227] ^ d[226] ^ d[225] ^ d[223] ^ d[221] ^ d[220] ^ d[219] ^ d[215] ^ d[214] ^ d[210] ^ d[207] ^ d[204] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[194] ^ d[192] ^ d[191] ^ d[190] ^ d[189] ^ d[187] ^ d[181] ^ d[180] ^ d[178] ^ d[175] ^ d[174] ^ d[173] ^ d[171] ^ d[169] ^ d[164] ^ d[161] ^ d[159] ^ d[153] ^ d[149] ^ d[147] ^ d[146] ^ d[145] ^ d[144] ^ d[142] ^ d[137] ^ d[135] ^ d[134] ^ d[127] ^ d[126] ^ d[125] ^ d[123] ^ d[122] ^ d[121] ^ d[118] ^ d[115] ^ d[113] ^ d[111] ^ d[109] ^ d[106] ^ d[105] ^ d[104] ^ d[103] ^ d[99] ^ d[98] ^ d[97] ^ d[86] ^ d[84] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[71] ^ d[70] ^ d[69] ^ d[65] ^ d[64] ^ d[62] ^ d[60] ^ d[58] ^ d[57] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[50] ^ d[49] ^ d[48] ^ d[46] ^ d[44] ^ d[43] ^ d[42] ^ d[41] ^ d[39] ^ d[38] ^ d[36] ^ d[32] ^ d[31] ^ d[30] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[15] ^ d[12] ^ d[10] ^ d[7] ^ d[6] ^ d[5] ^ d[2] ^ d[1] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[6] ^ c[7] ^ c[8] ^ c[10] ^ c[11] ^ c[14] ^ c[15] ^ c[17] ^ c[18] ^ c[20] ^ c[21];
    crc_func_0 = newcrc;
  end
  endfunction

////////////////////////////////////////////////////////////////////////////////
// Copyright (C) 1999-2008 Easics NV.
// This source file may be used and distributed without restriction
// provided that this copyright statement is not removed from the file
// and that any derivative work contains the original copyright notice
// and the associated disclaimer.
//
// THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
// WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
//
// Purpose : synthesizable CRC function
//   * polynomial: (0 1 3 4 5 6 7 10 11 14 17 18 23)
//   * data width: 256
//
// Info : tools@easics.be
//        http://www.easics.com
////////////////////////////////////////////////////////////////////////////////

  // polynomial: (0 1 3 4 5 6 7 10 11 14 17 18 23)
  // data width: 256
  // convention: the first serial bit is D[255]
  function [22:0] crc_func_1;

    input [255:0] Data;
    input [22:0] crc;
    reg [255:0] d;
    reg [22:0] c;
    reg [22:0] newcrc;
  begin
    d = Data;
    c = crc;

    newcrc[0] = d[255] ^ d[254] ^ d[252] ^ d[249] ^ d[248] ^ d[246] ^ d[245] ^ d[243] ^ d[242] ^ d[240] ^ d[239] ^ d[238] ^ d[236] ^ d[235] ^ d[232] ^ d[231] ^ d[230] ^ d[229] ^ d[228] ^ d[225] ^ d[223] ^ d[222] ^ d[219] ^ d[218] ^ d[217] ^ d[215] ^ d[213] ^ d[211] ^ d[210] ^ d[207] ^ d[206] ^ d[203] ^ d[195] ^ d[194] ^ d[193] ^ d[190] ^ d[189] ^ d[184] ^ d[178] ^ d[176] ^ d[172] ^ d[171] ^ d[168] ^ d[166] ^ d[165] ^ d[162] ^ d[158] ^ d[154] ^ d[152] ^ d[148] ^ d[147] ^ d[144] ^ d[143] ^ d[142] ^ d[140] ^ d[139] ^ d[137] ^ d[136] ^ d[133] ^ d[131] ^ d[129] ^ d[128] ^ d[127] ^ d[126] ^ d[125] ^ d[124] ^ d[122] ^ d[121] ^ d[119] ^ d[117] ^ d[115] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[109] ^ d[108] ^ d[107] ^ d[104] ^ d[103] ^ d[98] ^ d[96] ^ d[95] ^ d[94] ^ d[93] ^ d[92] ^ d[87] ^ d[86] ^ d[84] ^ d[83] ^ d[81] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[74] ^ d[72] ^ d[71] ^ d[68] ^ d[66] ^ d[65] ^ d[62] ^ d[60] ^ d[59] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[50] ^ d[49] ^ d[46] ^ d[44] ^ d[43] ^ d[42] ^ d[39] ^ d[38] ^ d[31] ^ d[29] ^ d[26] ^ d[23] ^ d[21] ^ d[18] ^ d[15] ^ d[13] ^ d[10] ^ d[9] ^ d[6] ^ d[5] ^ d[0] ^ c[2] ^ c[3] ^ c[5] ^ c[6] ^ c[7] ^ c[9] ^ c[10] ^ c[12] ^ c[13] ^ c[15] ^ c[16] ^ c[19] ^ c[21] ^ c[22];
    newcrc[1] = d[254] ^ d[253] ^ d[252] ^ d[250] ^ d[248] ^ d[247] ^ d[245] ^ d[244] ^ d[242] ^ d[241] ^ d[238] ^ d[237] ^ d[235] ^ d[233] ^ d[228] ^ d[226] ^ d[225] ^ d[224] ^ d[222] ^ d[220] ^ d[217] ^ d[216] ^ d[215] ^ d[214] ^ d[213] ^ d[212] ^ d[210] ^ d[208] ^ d[206] ^ d[204] ^ d[203] ^ d[196] ^ d[193] ^ d[191] ^ d[189] ^ d[185] ^ d[184] ^ d[179] ^ d[178] ^ d[177] ^ d[176] ^ d[173] ^ d[171] ^ d[169] ^ d[168] ^ d[167] ^ d[165] ^ d[163] ^ d[162] ^ d[159] ^ d[158] ^ d[155] ^ d[154] ^ d[153] ^ d[152] ^ d[149] ^ d[147] ^ d[145] ^ d[142] ^ d[141] ^ d[139] ^ d[138] ^ d[136] ^ d[134] ^ d[133] ^ d[132] ^ d[131] ^ d[130] ^ d[124] ^ d[123] ^ d[121] ^ d[120] ^ d[119] ^ d[118] ^ d[117] ^ d[116] ^ d[111] ^ d[110] ^ d[107] ^ d[105] ^ d[103] ^ d[99] ^ d[98] ^ d[97] ^ d[92] ^ d[88] ^ d[86] ^ d[85] ^ d[83] ^ d[82] ^ d[81] ^ d[80] ^ d[77] ^ d[76] ^ d[74] ^ d[73] ^ d[71] ^ d[69] ^ d[68] ^ d[67] ^ d[65] ^ d[63] ^ d[62] ^ d[61] ^ d[55] ^ d[51] ^ d[49] ^ d[47] ^ d[46] ^ d[45] ^ d[42] ^ d[40] ^ d[38] ^ d[32] ^ d[31] ^ d[30] ^ d[29] ^ d[27] ^ d[26] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[19] ^ d[18] ^ d[16] ^ d[15] ^ d[14] ^ d[13] ^ d[11] ^ d[9] ^ d[7] ^ d[5] ^ d[1] ^ d[0] ^ c[0] ^ c[2] ^ c[4] ^ c[5] ^ c[8] ^ c[9] ^ c[11] ^ c[12] ^ c[14] ^ c[15] ^ c[17] ^ c[19] ^ c[20] ^ c[21];
    newcrc[2] = d[255] ^ d[254] ^ d[253] ^ d[251] ^ d[249] ^ d[248] ^ d[246] ^ d[245] ^ d[243] ^ d[242] ^ d[239] ^ d[238] ^ d[236] ^ d[234] ^ d[229] ^ d[227] ^ d[226] ^ d[225] ^ d[223] ^ d[221] ^ d[218] ^ d[217] ^ d[216] ^ d[215] ^ d[214] ^ d[213] ^ d[211] ^ d[209] ^ d[207] ^ d[205] ^ d[204] ^ d[197] ^ d[194] ^ d[192] ^ d[190] ^ d[186] ^ d[185] ^ d[180] ^ d[179] ^ d[178] ^ d[177] ^ d[174] ^ d[172] ^ d[170] ^ d[169] ^ d[168] ^ d[166] ^ d[164] ^ d[163] ^ d[160] ^ d[159] ^ d[156] ^ d[155] ^ d[154] ^ d[153] ^ d[150] ^ d[148] ^ d[146] ^ d[143] ^ d[142] ^ d[140] ^ d[139] ^ d[137] ^ d[135] ^ d[134] ^ d[133] ^ d[132] ^ d[131] ^ d[125] ^ d[124] ^ d[122] ^ d[121] ^ d[120] ^ d[119] ^ d[118] ^ d[117] ^ d[112] ^ d[111] ^ d[108] ^ d[106] ^ d[104] ^ d[100] ^ d[99] ^ d[98] ^ d[93] ^ d[89] ^ d[87] ^ d[86] ^ d[84] ^ d[83] ^ d[82] ^ d[81] ^ d[78] ^ d[77] ^ d[75] ^ d[74] ^ d[72] ^ d[70] ^ d[69] ^ d[68] ^ d[66] ^ d[64] ^ d[63] ^ d[62] ^ d[56] ^ d[52] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[43] ^ d[41] ^ d[39] ^ d[33] ^ d[32] ^ d[31] ^ d[30] ^ d[28] ^ d[27] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[20] ^ d[19] ^ d[17] ^ d[16] ^ d[15] ^ d[14] ^ d[12] ^ d[10] ^ d[8] ^ d[6] ^ d[2] ^ d[1] ^ c[1] ^ c[3] ^ c[5] ^ c[6] ^ c[9] ^ c[10] ^ c[12] ^ c[13] ^ c[15] ^ c[16] ^ c[18] ^ c[20] ^ c[21] ^ c[22];
    newcrc[3] = d[250] ^ d[248] ^ d[247] ^ d[245] ^ d[244] ^ d[242] ^ d[238] ^ d[237] ^ d[236] ^ d[232] ^ d[231] ^ d[229] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[216] ^ d[214] ^ d[213] ^ d[212] ^ d[211] ^ d[208] ^ d[207] ^ d[205] ^ d[203] ^ d[198] ^ d[194] ^ d[191] ^ d[190] ^ d[189] ^ d[187] ^ d[186] ^ d[184] ^ d[181] ^ d[180] ^ d[179] ^ d[176] ^ d[175] ^ d[173] ^ d[172] ^ d[170] ^ d[169] ^ d[168] ^ d[167] ^ d[166] ^ d[164] ^ d[162] ^ d[161] ^ d[160] ^ d[158] ^ d[157] ^ d[156] ^ d[155] ^ d[152] ^ d[151] ^ d[149] ^ d[148] ^ d[142] ^ d[141] ^ d[139] ^ d[138] ^ d[137] ^ d[135] ^ d[134] ^ d[132] ^ d[131] ^ d[129] ^ d[128] ^ d[127] ^ d[124] ^ d[123] ^ d[120] ^ d[118] ^ d[117] ^ d[115] ^ d[114] ^ d[111] ^ d[108] ^ d[105] ^ d[104] ^ d[103] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[96] ^ d[95] ^ d[93] ^ d[92] ^ d[90] ^ d[88] ^ d[86] ^ d[85] ^ d[82] ^ d[81] ^ d[77] ^ d[76] ^ d[74] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[64] ^ d[63] ^ d[62] ^ d[60] ^ d[59] ^ d[58] ^ d[56] ^ d[55] ^ d[53] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[43] ^ d[40] ^ d[39] ^ d[38] ^ d[34] ^ d[33] ^ d[32] ^ d[28] ^ d[25] ^ d[24] ^ d[20] ^ d[17] ^ d[16] ^ d[11] ^ d[10] ^ d[7] ^ d[6] ^ d[5] ^ d[3] ^ d[2] ^ d[0] ^ c[3] ^ c[4] ^ c[5] ^ c[9] ^ c[11] ^ c[12] ^ c[14] ^ c[15] ^ c[17];
    newcrc[4] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[242] ^ d[240] ^ d[237] ^ d[236] ^ d[235] ^ d[233] ^ d[231] ^ d[229] ^ d[227] ^ d[226] ^ d[224] ^ d[223] ^ d[222] ^ d[219] ^ d[218] ^ d[214] ^ d[212] ^ d[211] ^ d[210] ^ d[209] ^ d[208] ^ d[207] ^ d[204] ^ d[203] ^ d[199] ^ d[194] ^ d[193] ^ d[192] ^ d[191] ^ d[189] ^ d[188] ^ d[187] ^ d[185] ^ d[184] ^ d[182] ^ d[181] ^ d[180] ^ d[178] ^ d[177] ^ d[174] ^ d[173] ^ d[172] ^ d[170] ^ d[169] ^ d[167] ^ d[166] ^ d[163] ^ d[161] ^ d[159] ^ d[157] ^ d[156] ^ d[154] ^ d[153] ^ d[150] ^ d[149] ^ d[148] ^ d[147] ^ d[144] ^ d[138] ^ d[137] ^ d[135] ^ d[132] ^ d[131] ^ d[130] ^ d[127] ^ d[126] ^ d[122] ^ d[118] ^ d[117] ^ d[116] ^ d[114] ^ d[113] ^ d[111] ^ d[108] ^ d[107] ^ d[106] ^ d[105] ^ d[103] ^ d[102] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[97] ^ d[95] ^ d[92] ^ d[91] ^ d[89] ^ d[84] ^ d[82] ^ d[81] ^ d[79] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[67] ^ d[66] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[58] ^ d[55] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[43] ^ d[42] ^ d[41] ^ d[40] ^ d[38] ^ d[35] ^ d[34] ^ d[33] ^ d[31] ^ d[25] ^ d[23] ^ d[17] ^ d[15] ^ d[13] ^ d[12] ^ d[11] ^ d[10] ^ d[9] ^ d[8] ^ d[7] ^ d[5] ^ d[4] ^ d[3] ^ d[1] ^ d[0] ^ c[0] ^ c[2] ^ c[3] ^ c[4] ^ c[7] ^ c[9] ^ c[18] ^ c[19] ^ c[21] ^ c[22];
    newcrc[5] = d[254] ^ d[253] ^ d[249] ^ d[248] ^ d[246] ^ d[245] ^ d[242] ^ d[241] ^ d[240] ^ d[239] ^ d[237] ^ d[235] ^ d[234] ^ d[231] ^ d[229] ^ d[227] ^ d[224] ^ d[222] ^ d[220] ^ d[218] ^ d[217] ^ d[212] ^ d[209] ^ d[208] ^ d[207] ^ d[206] ^ d[205] ^ d[204] ^ d[203] ^ d[200] ^ d[192] ^ d[188] ^ d[186] ^ d[185] ^ d[184] ^ d[183] ^ d[182] ^ d[181] ^ d[179] ^ d[176] ^ d[175] ^ d[174] ^ d[173] ^ d[172] ^ d[170] ^ d[167] ^ d[166] ^ d[165] ^ d[164] ^ d[160] ^ d[157] ^ d[155] ^ d[152] ^ d[151] ^ d[150] ^ d[149] ^ d[147] ^ d[145] ^ d[144] ^ d[143] ^ d[142] ^ d[140] ^ d[138] ^ d[137] ^ d[132] ^ d[129] ^ d[126] ^ d[125] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[118] ^ d[113] ^ d[111] ^ d[106] ^ d[102] ^ d[101] ^ d[100] ^ d[99] ^ d[95] ^ d[94] ^ d[90] ^ d[87] ^ d[86] ^ d[85] ^ d[84] ^ d[82] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[73] ^ d[72] ^ d[70] ^ d[67] ^ d[66] ^ d[64] ^ d[63] ^ d[60] ^ d[58] ^ d[57] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[41] ^ d[38] ^ d[36] ^ d[35] ^ d[34] ^ d[32] ^ d[31] ^ d[29] ^ d[24] ^ d[23] ^ d[21] ^ d[16] ^ d[15] ^ d[14] ^ d[12] ^ d[11] ^ d[8] ^ d[4] ^ d[2] ^ d[1] ^ d[0] ^ c[1] ^ c[2] ^ c[4] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[12] ^ c[13] ^ c[15] ^ c[16] ^ c[20] ^ c[21];
    newcrc[6] = d[252] ^ d[250] ^ d[248] ^ d[247] ^ d[245] ^ d[241] ^ d[239] ^ d[231] ^ d[229] ^ d[222] ^ d[221] ^ d[217] ^ d[215] ^ d[211] ^ d[209] ^ d[208] ^ d[205] ^ d[204] ^ d[203] ^ d[201] ^ d[195] ^ d[194] ^ d[190] ^ d[187] ^ d[186] ^ d[185] ^ d[183] ^ d[182] ^ d[180] ^ d[178] ^ d[177] ^ d[175] ^ d[174] ^ d[173] ^ d[172] ^ d[167] ^ d[162] ^ d[161] ^ d[156] ^ d[154] ^ d[153] ^ d[151] ^ d[150] ^ d[147] ^ d[146] ^ d[145] ^ d[142] ^ d[141] ^ d[140] ^ d[138] ^ d[137] ^ d[136] ^ d[131] ^ d[130] ^ d[129] ^ d[128] ^ d[123] ^ d[121] ^ d[117] ^ d[115] ^ d[113] ^ d[111] ^ d[109] ^ d[108] ^ d[104] ^ d[102] ^ d[101] ^ d[100] ^ d[98] ^ d[94] ^ d[93] ^ d[92] ^ d[91] ^ d[88] ^ d[85] ^ d[84] ^ d[82] ^ d[80] ^ d[77] ^ d[76] ^ d[75] ^ d[73] ^ d[72] ^ d[67] ^ d[66] ^ d[64] ^ d[62] ^ d[61] ^ d[60] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[44] ^ d[43] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[33] ^ d[32] ^ d[31] ^ d[30] ^ d[29] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[18] ^ d[17] ^ d[16] ^ d[12] ^ d[10] ^ d[6] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[6] ^ c[8] ^ c[12] ^ c[14] ^ c[15] ^ c[17] ^ c[19];
    newcrc[7] = d[255] ^ d[254] ^ d[253] ^ d[252] ^ d[251] ^ d[245] ^ d[243] ^ d[239] ^ d[238] ^ d[236] ^ d[235] ^ d[231] ^ d[229] ^ d[228] ^ d[225] ^ d[219] ^ d[217] ^ d[216] ^ d[215] ^ d[213] ^ d[212] ^ d[211] ^ d[209] ^ d[207] ^ d[205] ^ d[204] ^ d[203] ^ d[202] ^ d[196] ^ d[194] ^ d[193] ^ d[191] ^ d[190] ^ d[189] ^ d[188] ^ d[187] ^ d[186] ^ d[183] ^ d[181] ^ d[179] ^ d[175] ^ d[174] ^ d[173] ^ d[172] ^ d[171] ^ d[166] ^ d[165] ^ d[163] ^ d[158] ^ d[157] ^ d[155] ^ d[151] ^ d[146] ^ d[144] ^ d[141] ^ d[140] ^ d[138] ^ d[136] ^ d[133] ^ d[132] ^ d[130] ^ d[128] ^ d[127] ^ d[126] ^ d[125] ^ d[121] ^ d[119] ^ d[118] ^ d[117] ^ d[116] ^ d[115] ^ d[113] ^ d[111] ^ d[110] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[102] ^ d[101] ^ d[99] ^ d[98] ^ d[96] ^ d[89] ^ d[87] ^ d[85] ^ d[84] ^ d[79] ^ d[76] ^ d[75] ^ d[73] ^ d[72] ^ d[71] ^ d[67] ^ d[66] ^ d[63] ^ d[61] ^ d[60] ^ d[59] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[45] ^ d[43] ^ d[42] ^ d[37] ^ d[36] ^ d[34] ^ d[33] ^ d[32] ^ d[30] ^ d[29] ^ d[27] ^ d[25] ^ d[24] ^ d[22] ^ d[21] ^ d[19] ^ d[17] ^ d[15] ^ d[11] ^ d[10] ^ d[9] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[2] ^ c[3] ^ c[5] ^ c[6] ^ c[10] ^ c[12] ^ c[18] ^ c[19] ^ c[20] ^ c[21] ^ c[22];
    newcrc[8] = d[255] ^ d[254] ^ d[253] ^ d[252] ^ d[246] ^ d[244] ^ d[240] ^ d[239] ^ d[237] ^ d[236] ^ d[232] ^ d[230] ^ d[229] ^ d[226] ^ d[220] ^ d[218] ^ d[217] ^ d[216] ^ d[214] ^ d[213] ^ d[212] ^ d[210] ^ d[208] ^ d[206] ^ d[205] ^ d[204] ^ d[203] ^ d[197] ^ d[195] ^ d[194] ^ d[192] ^ d[191] ^ d[190] ^ d[189] ^ d[188] ^ d[187] ^ d[184] ^ d[182] ^ d[180] ^ d[176] ^ d[175] ^ d[174] ^ d[173] ^ d[172] ^ d[167] ^ d[166] ^ d[164] ^ d[159] ^ d[158] ^ d[156] ^ d[152] ^ d[147] ^ d[145] ^ d[142] ^ d[141] ^ d[139] ^ d[137] ^ d[134] ^ d[133] ^ d[131] ^ d[129] ^ d[128] ^ d[127] ^ d[126] ^ d[122] ^ d[120] ^ d[119] ^ d[118] ^ d[117] ^ d[116] ^ d[114] ^ d[112] ^ d[111] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[103] ^ d[102] ^ d[100] ^ d[99] ^ d[97] ^ d[90] ^ d[88] ^ d[86] ^ d[85] ^ d[80] ^ d[77] ^ d[76] ^ d[74] ^ d[73] ^ d[72] ^ d[68] ^ d[67] ^ d[64] ^ d[62] ^ d[61] ^ d[60] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[49] ^ d[48] ^ d[47] ^ d[46] ^ d[44] ^ d[43] ^ d[38] ^ d[37] ^ d[35] ^ d[34] ^ d[33] ^ d[31] ^ d[30] ^ d[28] ^ d[26] ^ d[25] ^ d[23] ^ d[22] ^ d[20] ^ d[18] ^ d[16] ^ d[12] ^ d[11] ^ d[10] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ c[3] ^ c[4] ^ c[6] ^ c[7] ^ c[11] ^ c[13] ^ c[19] ^ c[20] ^ c[21] ^ c[22];
    newcrc[9] = d[255] ^ d[254] ^ d[253] ^ d[247] ^ d[245] ^ d[241] ^ d[240] ^ d[238] ^ d[237] ^ d[233] ^ d[231] ^ d[230] ^ d[227] ^ d[221] ^ d[219] ^ d[218] ^ d[217] ^ d[215] ^ d[214] ^ d[213] ^ d[211] ^ d[209] ^ d[207] ^ d[206] ^ d[205] ^ d[204] ^ d[198] ^ d[196] ^ d[195] ^ d[193] ^ d[192] ^ d[191] ^ d[190] ^ d[189] ^ d[188] ^ d[185] ^ d[183] ^ d[181] ^ d[177] ^ d[176] ^ d[175] ^ d[174] ^ d[173] ^ d[168] ^ d[167] ^ d[165] ^ d[160] ^ d[159] ^ d[157] ^ d[153] ^ d[148] ^ d[146] ^ d[143] ^ d[142] ^ d[140] ^ d[138] ^ d[135] ^ d[134] ^ d[132] ^ d[130] ^ d[129] ^ d[128] ^ d[127] ^ d[123] ^ d[121] ^ d[120] ^ d[119] ^ d[118] ^ d[117] ^ d[115] ^ d[113] ^ d[112] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[104] ^ d[103] ^ d[101] ^ d[100] ^ d[98] ^ d[91] ^ d[89] ^ d[87] ^ d[86] ^ d[81] ^ d[78] ^ d[77] ^ d[75] ^ d[74] ^ d[73] ^ d[69] ^ d[68] ^ d[65] ^ d[63] ^ d[62] ^ d[61] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[50] ^ d[49] ^ d[48] ^ d[47] ^ d[45] ^ d[44] ^ d[39] ^ d[38] ^ d[36] ^ d[35] ^ d[34] ^ d[32] ^ d[31] ^ d[29] ^ d[27] ^ d[26] ^ d[24] ^ d[23] ^ d[21] ^ d[19] ^ d[17] ^ d[13] ^ d[12] ^ d[11] ^ d[9] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ c[0] ^ c[4] ^ c[5] ^ c[7] ^ c[8] ^ c[12] ^ c[14] ^ c[20] ^ c[21] ^ c[22];
    newcrc[10] = d[252] ^ d[249] ^ d[245] ^ d[243] ^ d[241] ^ d[240] ^ d[236] ^ d[235] ^ d[234] ^ d[230] ^ d[229] ^ d[225] ^ d[223] ^ d[220] ^ d[217] ^ d[216] ^ d[214] ^ d[213] ^ d[212] ^ d[211] ^ d[208] ^ d[205] ^ d[203] ^ d[199] ^ d[197] ^ d[196] ^ d[195] ^ d[192] ^ d[191] ^ d[186] ^ d[182] ^ d[177] ^ d[175] ^ d[174] ^ d[172] ^ d[171] ^ d[169] ^ d[165] ^ d[162] ^ d[161] ^ d[160] ^ d[152] ^ d[149] ^ d[148] ^ d[142] ^ d[141] ^ d[140] ^ d[137] ^ d[135] ^ d[130] ^ d[127] ^ d[126] ^ d[125] ^ d[120] ^ d[118] ^ d[117] ^ d[116] ^ d[115] ^ d[112] ^ d[110] ^ d[109] ^ d[105] ^ d[103] ^ d[102] ^ d[101] ^ d[99] ^ d[98] ^ d[96] ^ d[95] ^ d[94] ^ d[93] ^ d[90] ^ d[88] ^ d[86] ^ d[84] ^ d[83] ^ d[82] ^ d[81] ^ d[77] ^ d[76] ^ d[72] ^ d[71] ^ d[70] ^ d[69] ^ d[68] ^ d[65] ^ d[64] ^ d[63] ^ d[60] ^ d[59] ^ d[58] ^ d[54] ^ d[53] ^ d[51] ^ d[48] ^ d[45] ^ d[44] ^ d[43] ^ d[42] ^ d[40] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[33] ^ d[32] ^ d[31] ^ d[30] ^ d[29] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[15] ^ d[14] ^ d[12] ^ d[8] ^ d[7] ^ d[4] ^ d[3] ^ d[0] ^ c[1] ^ c[2] ^ c[3] ^ c[7] ^ c[8] ^ c[10] ^ c[12] ^ c[16] ^ c[19];
    newcrc[11] = d[255] ^ d[254] ^ d[253] ^ d[252] ^ d[250] ^ d[249] ^ d[248] ^ d[245] ^ d[244] ^ d[243] ^ d[241] ^ d[240] ^ d[239] ^ d[238] ^ d[237] ^ d[232] ^ d[229] ^ d[228] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[222] ^ d[221] ^ d[219] ^ d[214] ^ d[212] ^ d[211] ^ d[210] ^ d[209] ^ d[207] ^ d[204] ^ d[203] ^ d[200] ^ d[198] ^ d[197] ^ d[196] ^ d[195] ^ d[194] ^ d[192] ^ d[190] ^ d[189] ^ d[187] ^ d[184] ^ d[183] ^ d[175] ^ d[173] ^ d[171] ^ d[170] ^ d[168] ^ d[165] ^ d[163] ^ d[161] ^ d[158] ^ d[154] ^ d[153] ^ d[152] ^ d[150] ^ d[149] ^ d[148] ^ d[147] ^ d[144] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[133] ^ d[129] ^ d[125] ^ d[124] ^ d[122] ^ d[118] ^ d[116] ^ d[115] ^ d[114] ^ d[112] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[102] ^ d[100] ^ d[99] ^ d[98] ^ d[97] ^ d[93] ^ d[92] ^ d[91] ^ d[89] ^ d[86] ^ d[85] ^ d[82] ^ d[81] ^ d[79] ^ d[75] ^ d[74] ^ d[73] ^ d[70] ^ d[69] ^ d[68] ^ d[64] ^ d[62] ^ d[61] ^ d[58] ^ d[57] ^ d[56] ^ d[54] ^ d[52] ^ d[50] ^ d[45] ^ d[42] ^ d[41] ^ d[37] ^ d[36] ^ d[34] ^ d[33] ^ d[32] ^ d[30] ^ d[28] ^ d[27] ^ d[25] ^ d[24] ^ d[22] ^ d[18] ^ d[16] ^ d[10] ^ d[8] ^ d[6] ^ d[4] ^ d[1] ^ d[0] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[10] ^ c[11] ^ c[12] ^ c[15] ^ c[16] ^ c[17] ^ c[19] ^ c[20] ^ c[21] ^ c[22];
    newcrc[12] = d[255] ^ d[254] ^ d[253] ^ d[251] ^ d[250] ^ d[249] ^ d[246] ^ d[245] ^ d[244] ^ d[242] ^ d[241] ^ d[240] ^ d[239] ^ d[238] ^ d[233] ^ d[230] ^ d[229] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[222] ^ d[220] ^ d[215] ^ d[213] ^ d[212] ^ d[211] ^ d[210] ^ d[208] ^ d[205] ^ d[204] ^ d[201] ^ d[199] ^ d[198] ^ d[197] ^ d[196] ^ d[195] ^ d[193] ^ d[191] ^ d[190] ^ d[188] ^ d[185] ^ d[184] ^ d[176] ^ d[174] ^ d[172] ^ d[171] ^ d[169] ^ d[166] ^ d[164] ^ d[162] ^ d[159] ^ d[155] ^ d[154] ^ d[153] ^ d[151] ^ d[150] ^ d[149] ^ d[148] ^ d[145] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[134] ^ d[130] ^ d[126] ^ d[125] ^ d[123] ^ d[119] ^ d[117] ^ d[116] ^ d[115] ^ d[113] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[103] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[94] ^ d[93] ^ d[92] ^ d[90] ^ d[87] ^ d[86] ^ d[83] ^ d[82] ^ d[80] ^ d[76] ^ d[75] ^ d[74] ^ d[71] ^ d[70] ^ d[69] ^ d[65] ^ d[63] ^ d[62] ^ d[59] ^ d[58] ^ d[57] ^ d[55] ^ d[53] ^ d[51] ^ d[46] ^ d[43] ^ d[42] ^ d[38] ^ d[37] ^ d[35] ^ d[34] ^ d[33] ^ d[31] ^ d[29] ^ d[28] ^ d[26] ^ d[25] ^ d[23] ^ d[19] ^ d[17] ^ d[11] ^ d[9] ^ d[7] ^ d[5] ^ d[2] ^ d[1] ^ c[0] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[11] ^ c[12] ^ c[13] ^ c[16] ^ c[17] ^ c[18] ^ c[20] ^ c[21] ^ c[22];
    newcrc[13] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[250] ^ d[247] ^ d[246] ^ d[245] ^ d[243] ^ d[242] ^ d[241] ^ d[240] ^ d[239] ^ d[234] ^ d[231] ^ d[230] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[221] ^ d[216] ^ d[214] ^ d[213] ^ d[212] ^ d[211] ^ d[209] ^ d[206] ^ d[205] ^ d[202] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[196] ^ d[194] ^ d[192] ^ d[191] ^ d[189] ^ d[186] ^ d[185] ^ d[177] ^ d[175] ^ d[173] ^ d[172] ^ d[170] ^ d[167] ^ d[165] ^ d[163] ^ d[160] ^ d[156] ^ d[155] ^ d[154] ^ d[152] ^ d[151] ^ d[150] ^ d[149] ^ d[146] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[135] ^ d[131] ^ d[127] ^ d[126] ^ d[124] ^ d[120] ^ d[118] ^ d[117] ^ d[116] ^ d[114] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[104] ^ d[102] ^ d[101] ^ d[100] ^ d[99] ^ d[95] ^ d[94] ^ d[93] ^ d[91] ^ d[88] ^ d[87] ^ d[84] ^ d[83] ^ d[81] ^ d[77] ^ d[76] ^ d[75] ^ d[72] ^ d[71] ^ d[70] ^ d[66] ^ d[64] ^ d[63] ^ d[60] ^ d[59] ^ d[58] ^ d[56] ^ d[54] ^ d[52] ^ d[47] ^ d[44] ^ d[43] ^ d[39] ^ d[38] ^ d[36] ^ d[35] ^ d[34] ^ d[32] ^ d[30] ^ d[29] ^ d[27] ^ d[26] ^ d[24] ^ d[20] ^ d[18] ^ d[12] ^ d[10] ^ d[8] ^ d[6] ^ d[3] ^ d[2] ^ c[1] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[12] ^ c[13] ^ c[14] ^ c[17] ^ c[18] ^ c[19] ^ c[21] ^ c[22];
    newcrc[14] = d[254] ^ d[253] ^ d[251] ^ d[249] ^ d[247] ^ d[245] ^ d[244] ^ d[241] ^ d[239] ^ d[238] ^ d[236] ^ d[230] ^ d[227] ^ d[226] ^ d[224] ^ d[223] ^ d[219] ^ d[218] ^ d[214] ^ d[212] ^ d[211] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[194] ^ d[192] ^ d[189] ^ d[187] ^ d[186] ^ d[184] ^ d[174] ^ d[173] ^ d[172] ^ d[165] ^ d[164] ^ d[162] ^ d[161] ^ d[158] ^ d[157] ^ d[156] ^ d[155] ^ d[154] ^ d[153] ^ d[151] ^ d[150] ^ d[148] ^ d[141] ^ d[139] ^ d[137] ^ d[133] ^ d[132] ^ d[131] ^ d[129] ^ d[126] ^ d[124] ^ d[122] ^ d[118] ^ d[114] ^ d[110] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[102] ^ d[101] ^ d[100] ^ d[98] ^ d[93] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[85] ^ d[83] ^ d[82] ^ d[81] ^ d[79] ^ d[76] ^ d[75] ^ d[74] ^ d[73] ^ d[68] ^ d[67] ^ d[66] ^ d[64] ^ d[62] ^ d[61] ^ d[58] ^ d[56] ^ d[53] ^ d[50] ^ d[49] ^ d[48] ^ d[46] ^ d[45] ^ d[43] ^ d[42] ^ d[40] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[33] ^ d[30] ^ d[29] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[23] ^ d[19] ^ d[18] ^ d[15] ^ d[11] ^ d[10] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[0] ^ c[3] ^ c[5] ^ c[6] ^ c[8] ^ c[11] ^ c[12] ^ c[14] ^ c[16] ^ c[18] ^ c[20] ^ c[21];
    newcrc[15] = d[255] ^ d[254] ^ d[252] ^ d[250] ^ d[248] ^ d[246] ^ d[245] ^ d[242] ^ d[240] ^ d[239] ^ d[237] ^ d[231] ^ d[228] ^ d[227] ^ d[225] ^ d[224] ^ d[220] ^ d[219] ^ d[215] ^ d[213] ^ d[212] ^ d[202] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[195] ^ d[193] ^ d[190] ^ d[188] ^ d[187] ^ d[185] ^ d[175] ^ d[174] ^ d[173] ^ d[166] ^ d[165] ^ d[163] ^ d[162] ^ d[159] ^ d[158] ^ d[157] ^ d[156] ^ d[155] ^ d[154] ^ d[152] ^ d[151] ^ d[149] ^ d[142] ^ d[140] ^ d[138] ^ d[134] ^ d[133] ^ d[132] ^ d[130] ^ d[127] ^ d[125] ^ d[123] ^ d[119] ^ d[115] ^ d[111] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[103] ^ d[102] ^ d[101] ^ d[99] ^ d[94] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[84] ^ d[83] ^ d[82] ^ d[80] ^ d[77] ^ d[76] ^ d[75] ^ d[74] ^ d[69] ^ d[68] ^ d[67] ^ d[65] ^ d[63] ^ d[62] ^ d[59] ^ d[57] ^ d[54] ^ d[51] ^ d[50] ^ d[49] ^ d[47] ^ d[46] ^ d[44] ^ d[43] ^ d[41] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[34] ^ d[31] ^ d[30] ^ d[29] ^ d[28] ^ d[27] ^ d[26] ^ d[24] ^ d[20] ^ d[19] ^ d[16] ^ d[12] ^ d[11] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[1] ^ c[4] ^ c[6] ^ c[7] ^ c[9] ^ c[12] ^ c[13] ^ c[15] ^ c[17] ^ c[19] ^ c[21] ^ c[22];
    newcrc[16] = d[255] ^ d[253] ^ d[251] ^ d[249] ^ d[247] ^ d[246] ^ d[243] ^ d[241] ^ d[240] ^ d[238] ^ d[232] ^ d[229] ^ d[228] ^ d[226] ^ d[225] ^ d[221] ^ d[220] ^ d[216] ^ d[214] ^ d[213] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[199] ^ d[196] ^ d[194] ^ d[191] ^ d[189] ^ d[188] ^ d[186] ^ d[176] ^ d[175] ^ d[174] ^ d[167] ^ d[166] ^ d[164] ^ d[163] ^ d[160] ^ d[159] ^ d[158] ^ d[157] ^ d[156] ^ d[155] ^ d[153] ^ d[152] ^ d[150] ^ d[143] ^ d[141] ^ d[139] ^ d[135] ^ d[134] ^ d[133] ^ d[131] ^ d[128] ^ d[126] ^ d[124] ^ d[120] ^ d[116] ^ d[112] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[104] ^ d[103] ^ d[102] ^ d[100] ^ d[95] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[85] ^ d[84] ^ d[83] ^ d[81] ^ d[78] ^ d[77] ^ d[76] ^ d[75] ^ d[70] ^ d[69] ^ d[68] ^ d[66] ^ d[64] ^ d[63] ^ d[60] ^ d[58] ^ d[55] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[45] ^ d[44] ^ d[42] ^ d[40] ^ d[39] ^ d[38] ^ d[37] ^ d[35] ^ d[32] ^ d[31] ^ d[30] ^ d[29] ^ d[28] ^ d[27] ^ d[25] ^ d[21] ^ d[20] ^ d[17] ^ d[13] ^ d[12] ^ d[9] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[2] ^ c[5] ^ c[7] ^ c[8] ^ c[10] ^ c[13] ^ c[14] ^ c[16] ^ c[18] ^ c[20] ^ c[22];
    newcrc[17] = d[255] ^ d[250] ^ d[249] ^ d[247] ^ d[246] ^ d[245] ^ d[244] ^ d[243] ^ d[241] ^ d[240] ^ d[238] ^ d[236] ^ d[235] ^ d[233] ^ d[232] ^ d[231] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[223] ^ d[221] ^ d[219] ^ d[218] ^ d[214] ^ d[213] ^ d[211] ^ d[210] ^ d[207] ^ d[206] ^ d[204] ^ d[202] ^ d[201] ^ d[200] ^ d[197] ^ d[194] ^ d[193] ^ d[192] ^ d[187] ^ d[184] ^ d[178] ^ d[177] ^ d[175] ^ d[172] ^ d[171] ^ d[167] ^ d[166] ^ d[164] ^ d[162] ^ d[161] ^ d[160] ^ d[159] ^ d[157] ^ d[156] ^ d[153] ^ d[152] ^ d[151] ^ d[148] ^ d[147] ^ d[143] ^ d[139] ^ d[137] ^ d[135] ^ d[134] ^ d[133] ^ d[132] ^ d[131] ^ d[128] ^ d[126] ^ d[124] ^ d[122] ^ d[119] ^ d[115] ^ d[114] ^ d[112] ^ d[110] ^ d[109] ^ d[105] ^ d[101] ^ d[98] ^ d[95] ^ d[94] ^ d[93] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[85] ^ d[83] ^ d[82] ^ d[81] ^ d[76] ^ d[75] ^ d[74] ^ d[72] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[64] ^ d[62] ^ d[61] ^ d[60] ^ d[58] ^ d[57] ^ d[55] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[45] ^ d[44] ^ d[42] ^ d[41] ^ d[40] ^ d[36] ^ d[33] ^ d[32] ^ d[30] ^ d[28] ^ d[23] ^ d[22] ^ d[15] ^ d[14] ^ d[8] ^ d[7] ^ d[5] ^ d[3] ^ d[0] ^ c[0] ^ c[2] ^ c[3] ^ c[5] ^ c[7] ^ c[8] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[16] ^ c[17] ^ c[22];
    newcrc[18] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[250] ^ d[249] ^ d[247] ^ d[244] ^ d[243] ^ d[241] ^ d[240] ^ d[238] ^ d[237] ^ d[235] ^ d[234] ^ d[233] ^ d[231] ^ d[230] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[220] ^ d[218] ^ d[217] ^ d[214] ^ d[213] ^ d[212] ^ d[210] ^ d[208] ^ d[206] ^ d[205] ^ d[202] ^ d[201] ^ d[198] ^ d[190] ^ d[189] ^ d[188] ^ d[185] ^ d[184] ^ d[179] ^ d[173] ^ d[171] ^ d[167] ^ d[166] ^ d[163] ^ d[161] ^ d[160] ^ d[157] ^ d[153] ^ d[149] ^ d[147] ^ d[143] ^ d[142] ^ d[139] ^ d[138] ^ d[137] ^ d[135] ^ d[134] ^ d[132] ^ d[131] ^ d[128] ^ d[126] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[120] ^ d[119] ^ d[117] ^ d[116] ^ d[114] ^ d[112] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[104] ^ d[103] ^ d[102] ^ d[99] ^ d[98] ^ d[93] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[82] ^ d[81] ^ d[79] ^ d[78] ^ d[76] ^ d[74] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[67] ^ d[66] ^ d[63] ^ d[61] ^ d[60] ^ d[57] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[45] ^ d[44] ^ d[41] ^ d[39] ^ d[38] ^ d[37] ^ d[34] ^ d[33] ^ d[26] ^ d[24] ^ d[21] ^ d[18] ^ d[16] ^ d[13] ^ d[10] ^ d[8] ^ d[5] ^ d[4] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[4] ^ c[5] ^ c[7] ^ c[8] ^ c[10] ^ c[11] ^ c[14] ^ c[16] ^ c[17] ^ c[18] ^ c[19] ^ c[21] ^ c[22];
    newcrc[19] = d[255] ^ d[253] ^ d[252] ^ d[251] ^ d[250] ^ d[248] ^ d[245] ^ d[244] ^ d[242] ^ d[241] ^ d[239] ^ d[238] ^ d[236] ^ d[235] ^ d[234] ^ d[232] ^ d[231] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[221] ^ d[219] ^ d[218] ^ d[215] ^ d[214] ^ d[213] ^ d[211] ^ d[209] ^ d[207] ^ d[206] ^ d[203] ^ d[202] ^ d[199] ^ d[191] ^ d[190] ^ d[189] ^ d[186] ^ d[185] ^ d[180] ^ d[174] ^ d[172] ^ d[168] ^ d[167] ^ d[164] ^ d[162] ^ d[161] ^ d[158] ^ d[154] ^ d[150] ^ d[148] ^ d[144] ^ d[143] ^ d[140] ^ d[139] ^ d[138] ^ d[136] ^ d[135] ^ d[133] ^ d[132] ^ d[129] ^ d[127] ^ d[125] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[120] ^ d[118] ^ d[117] ^ d[115] ^ d[113] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[103] ^ d[100] ^ d[99] ^ d[94] ^ d[92] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[83] ^ d[82] ^ d[80] ^ d[79] ^ d[77] ^ d[75] ^ d[74] ^ d[73] ^ d[71] ^ d[70] ^ d[68] ^ d[67] ^ d[64] ^ d[62] ^ d[61] ^ d[58] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[46] ^ d[45] ^ d[42] ^ d[40] ^ d[39] ^ d[38] ^ d[35] ^ d[34] ^ d[27] ^ d[25] ^ d[22] ^ d[19] ^ d[17] ^ d[14] ^ d[11] ^ d[9] ^ d[6] ^ d[5] ^ d[2] ^ d[1] ^ c[1] ^ c[2] ^ c[3] ^ c[5] ^ c[6] ^ c[8] ^ c[9] ^ c[11] ^ c[12] ^ c[15] ^ c[17] ^ c[18] ^ c[19] ^ c[20] ^ c[22];
    newcrc[20] = d[254] ^ d[253] ^ d[252] ^ d[251] ^ d[249] ^ d[246] ^ d[245] ^ d[243] ^ d[242] ^ d[240] ^ d[239] ^ d[237] ^ d[236] ^ d[235] ^ d[233] ^ d[232] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[222] ^ d[220] ^ d[219] ^ d[216] ^ d[215] ^ d[214] ^ d[212] ^ d[210] ^ d[208] ^ d[207] ^ d[204] ^ d[203] ^ d[200] ^ d[192] ^ d[191] ^ d[190] ^ d[187] ^ d[186] ^ d[181] ^ d[175] ^ d[173] ^ d[169] ^ d[168] ^ d[165] ^ d[163] ^ d[162] ^ d[159] ^ d[155] ^ d[151] ^ d[149] ^ d[145] ^ d[144] ^ d[141] ^ d[140] ^ d[139] ^ d[137] ^ d[136] ^ d[134] ^ d[133] ^ d[130] ^ d[128] ^ d[126] ^ d[125] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[119] ^ d[118] ^ d[116] ^ d[114] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[104] ^ d[101] ^ d[100] ^ d[95] ^ d[93] ^ d[92] ^ d[91] ^ d[90] ^ d[89] ^ d[84] ^ d[83] ^ d[81] ^ d[80] ^ d[78] ^ d[76] ^ d[75] ^ d[74] ^ d[72] ^ d[71] ^ d[69] ^ d[68] ^ d[65] ^ d[63] ^ d[62] ^ d[59] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[47] ^ d[46] ^ d[43] ^ d[41] ^ d[40] ^ d[39] ^ d[36] ^ d[35] ^ d[28] ^ d[26] ^ d[23] ^ d[20] ^ d[18] ^ d[15] ^ d[12] ^ d[10] ^ d[7] ^ d[6] ^ d[3] ^ d[2] ^ c[0] ^ c[2] ^ c[3] ^ c[4] ^ c[6] ^ c[7] ^ c[9] ^ c[10] ^ c[12] ^ c[13] ^ c[16] ^ c[18] ^ c[19] ^ c[20] ^ c[21];
    newcrc[21] = d[255] ^ d[254] ^ d[253] ^ d[252] ^ d[250] ^ d[247] ^ d[246] ^ d[244] ^ d[243] ^ d[241] ^ d[240] ^ d[238] ^ d[237] ^ d[236] ^ d[234] ^ d[233] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[223] ^ d[221] ^ d[220] ^ d[217] ^ d[216] ^ d[215] ^ d[213] ^ d[211] ^ d[209] ^ d[208] ^ d[205] ^ d[204] ^ d[201] ^ d[193] ^ d[192] ^ d[191] ^ d[188] ^ d[187] ^ d[182] ^ d[176] ^ d[174] ^ d[170] ^ d[169] ^ d[166] ^ d[164] ^ d[163] ^ d[160] ^ d[156] ^ d[152] ^ d[150] ^ d[146] ^ d[145] ^ d[142] ^ d[141] ^ d[140] ^ d[138] ^ d[137] ^ d[135] ^ d[134] ^ d[131] ^ d[129] ^ d[127] ^ d[126] ^ d[125] ^ d[124] ^ d[123] ^ d[122] ^ d[120] ^ d[119] ^ d[117] ^ d[115] ^ d[113] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[105] ^ d[102] ^ d[101] ^ d[96] ^ d[94] ^ d[93] ^ d[92] ^ d[91] ^ d[90] ^ d[85] ^ d[84] ^ d[82] ^ d[81] ^ d[79] ^ d[77] ^ d[76] ^ d[75] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[66] ^ d[64] ^ d[63] ^ d[60] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[48] ^ d[47] ^ d[44] ^ d[42] ^ d[41] ^ d[40] ^ d[37] ^ d[36] ^ d[29] ^ d[27] ^ d[24] ^ d[21] ^ d[19] ^ d[16] ^ d[13] ^ d[11] ^ d[8] ^ d[7] ^ d[4] ^ d[3] ^ c[0] ^ c[1] ^ c[3] ^ c[4] ^ c[5] ^ c[7] ^ c[8] ^ c[10] ^ c[11] ^ c[13] ^ c[14] ^ c[17] ^ c[19] ^ c[20] ^ c[21] ^ c[22];
    newcrc[22] = d[255] ^ d[254] ^ d[253] ^ d[251] ^ d[248] ^ d[247] ^ d[245] ^ d[244] ^ d[242] ^ d[241] ^ d[239] ^ d[238] ^ d[237] ^ d[235] ^ d[234] ^ d[231] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[224] ^ d[222] ^ d[221] ^ d[218] ^ d[217] ^ d[216] ^ d[214] ^ d[212] ^ d[210] ^ d[209] ^ d[206] ^ d[205] ^ d[202] ^ d[194] ^ d[193] ^ d[192] ^ d[189] ^ d[188] ^ d[183] ^ d[177] ^ d[175] ^ d[171] ^ d[170] ^ d[167] ^ d[165] ^ d[164] ^ d[161] ^ d[157] ^ d[153] ^ d[151] ^ d[147] ^ d[146] ^ d[143] ^ d[142] ^ d[141] ^ d[139] ^ d[138] ^ d[136] ^ d[135] ^ d[132] ^ d[130] ^ d[128] ^ d[127] ^ d[126] ^ d[125] ^ d[124] ^ d[123] ^ d[121] ^ d[120] ^ d[118] ^ d[116] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[110] ^ d[108] ^ d[107] ^ d[106] ^ d[103] ^ d[102] ^ d[97] ^ d[95] ^ d[94] ^ d[93] ^ d[92] ^ d[91] ^ d[86] ^ d[85] ^ d[83] ^ d[82] ^ d[80] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[73] ^ d[71] ^ d[70] ^ d[67] ^ d[65] ^ d[64] ^ d[61] ^ d[59] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[49] ^ d[48] ^ d[45] ^ d[43] ^ d[42] ^ d[41] ^ d[38] ^ d[37] ^ d[30] ^ d[28] ^ d[25] ^ d[22] ^ d[20] ^ d[17] ^ d[14] ^ d[12] ^ d[9] ^ d[8] ^ d[5] ^ d[4] ^ c[1] ^ c[2] ^ c[4] ^ c[5] ^ c[6] ^ c[8] ^ c[9] ^ c[11] ^ c[12] ^ c[14] ^ c[15] ^ c[18] ^ c[20] ^ c[21] ^ c[22];
    crc_func_1 = newcrc;
  end
  endfunction


   wire [255:0] data_rev;
   wire [255:0] data_padded = {{(256-INPUT_WIDTH){1'b0}}, data};

   generate
      genvar 	i;
      for (i=0; i<32; i=i+1) begin: test
	 		assign data_rev[(31-i)*8 + 7 : (31-i)*8] = data_padded[i*8 + 7 : i*8];
      end
   endgenerate

   always @(posedge clk) begin
      if(reset) begin
	 		hash_0        <= 0;
	 		hash_1        <= 0;
      end else begin
	 		hash_0        <= crc_func_0(data_rev, 256'h0);
	 		hash_1        <= crc_func_1(data_rev, 256'h0);
      end // else: !if(reset)
   end
endmodule // hash
